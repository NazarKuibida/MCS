library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity transition_logic_int is

 Port ( CUR_STATE : in  std_logic_vector(2 downto 0);
           MODE : in  std_logic;
           RESET : in std_logic;
           NEXT_STATE : out  std_logic_vector(2 downto 0)
        );
		
end transition_logic_int;

architecture transition_logic_arc of transition_logic_int is

begin
    
NEXT_STATE(0) <=
    (not(RESET) and not(MODE) and not(CUR_STATE(2)) and not(CUR_STATE(1)) and not(CUR_STATE(0))) or
	 (not(RESET) and not(MODE) and not(CUR_STATE(2)) and CUR_STATE(1) and not(CUR_STATE(0))) or
	 (not(RESET) and not(MODE) and CUR_STATE(2) and not(CUR_STATE(1)) and not(CUR_STATE(0))) or
	 (not(RESET) and not(MODE) and CUR_STATE(2) and CUR_STATE(1) and not(CUR_STATE(0))) or
	 
	 (not(RESET) and MODE and CUR_STATE(2) and CUR_STATE(1) and not(CUR_STATE(0))) or
	 (not(RESET) and MODE and CUR_STATE(2) and not(CUR_STATE(1)) and not(CUR_STATE(0))) or
	 (not(RESET) and MODE and not(CUR_STATE(2)) and CUR_STATE(1) and not(CUR_STATE(0))) or
	 (not (RESET) and MODE and not(CUR_STATE(2)) and not(CUR_STATE(1)) and not(CUR_STATE(0)));
	 
	 
NEXT_STATE(1)<=
	 (not(RESET) and not(MODE) and not(CUR_STATE(2)) and not(CUR_STATE(1)) and CUR_STATE(0)) or
	 (not(RESET) and not(MODE) and not(CUR_STATE(2)) and CUR_STATE(1) and not(CUR_STATE(0))) or
	 (not(RESET) and not(MODE) and CUR_STATE(2) and not(CUR_STATE(1)) and CUR_STATE(0)) or
	 (not(RESET) and not(MODE) and CUR_STATE(2) and CUR_STATE(1) and not(CUR_STATE(0))) or
	 
	 
	 (not(RESET) and MODE and CUR_STATE(2) and CUR_STATE(1) and CUR_STATE(0)) or
	 (not(RESET) and MODE and CUR_STATE(2) and not(CUR_STATE(1)) and not(CUR_STATE(0))) or
	 (not(RESET) and MODE and not(CUR_STATE(2)) and CUR_STATE(1) and CUR_STATE(0)) or
	 (not (RESET) and MODE and not(CUR_STATE(2)) and not(CUR_STATE(1)) and not(CUR_STATE(0)));
	 
NEXT_STATE(2)<=
	 (not(RESET) and not(MODE) and not(CUR_STATE(2)) and CUR_STATE(1) and CUR_STATE(0)) or
	 (not(RESET) and not(MODE) and CUR_STATE(2) and not(CUR_STATE(1)) and not(CUR_STATE(0))) or
	 (not(RESET) and not(MODE) and CUR_STATE(2) and not(CUR_STATE(1)) and CUR_STATE(0)) or
	 (not(RESET) and not(MODE) and CUR_STATE(2) and CUR_STATE(1) and not(CUR_STATE(0))) or
	 
	 (not(RESET) and MODE and CUR_STATE(2) and CUR_STATE(1) and CUR_STATE(0)) or
	 (not(RESET) and MODE and CUR_STATE(2) and CUR_STATE(1) and not(CUR_STATE(0))) or
	 (not(RESET) and MODE and CUR_STATE(2) and not(CUR_STATE(1)) and CUR_STATE(0)) or
	 (not (RESET) and MODE and not(CUR_STATE(2)) and not(CUR_STATE(1)) and not(CUR_STATE(0)));
	 
             
end transition_logic_arc;




